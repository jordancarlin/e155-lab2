// lab2_tb.sv
// Jordan Carlin, jcarlin@hmc.edu, 7 September 2024
// Testbench for the E155 Lab 2 FPGA design

`timescale 1ns/1ns
`default_nettype none
`define N_TV 10

module lab2_tb();
  // Set up test signals
  logic        clk;
  logic [3:0]  s0, s1;
  logic [4:0]  leds;
  logic [6:0]  segs;
  logic        disp0, disp1;

  // Instantiate the device under test
  top dut(.*);

  // Generate clock signal with a period of 10 timesteps.
  always begin
    clk = 1; #5;
    clk = 0; #5;
  end


  // Apply test vectors
  initial begin
    #12;
    s0=4'b0000; s1=4'b0000; #20;
    s0=4'b0001; s1=4'b0000; #20;
    s0=4'b0000; s1=4'b0001; #20;
    s0=4'b0001; s1=4'b0001; #20;
    s0=4'b1111; s1=4'b0000; #20;
    s0=4'b0000; s1=4'b1111; #20;
    s0=4'b1111; s1=4'b1111; #20;
    s0=4'b0100; s1=4'b0010; #20;
  end

endmodule
